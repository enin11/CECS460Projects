`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:03:36 03/06/2018 
// Design Name: 
// Module Name:    TxRdy_Reg 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module TxRdy_Reg(input clk, rst
    output reg TxRdy);
	 
	 
	 	always @ (posedge clk, posedge rst)
		begin
			if (rst) 
				TxRdy <= 1'b1; else
			
			if (load == 1'b1 && done == 1'b1)
				TxRdy <= TxRdy; else
			
			if (done)
				TxRdy <= 1'b1; else
			
			if (load)
				TxRdy <= 1'b0;
			
			else
				TxRdy <= TxRdy; //for clarity
		end


endmodule
